----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    00:45:33 06/30/2020 
-- Design Name: 
-- Module Name:    register - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity register is
    Port ( clk : in  STD_LOGIC;
           rst : in  STD_LOGIC;
           regWrite : in  STD_LOGIC;
           Ra : in  STD_LOGIC_VECTOR (2 downto 0);
           Rb : in  STD_LOGIC_VECTOR (2 downto 0);
           Rw : in  STD_LOGIC_VECTOR (2 downto 0);
           din : in  STD_LOGIC_VECTOR (15 downto 0);
           doutA : out  STD_LOGIC_VECTOR (15 downto 0);
           doutB : out  STD_LOGIC_VECTOR (15 downto 0));
end register;

architecture Behavioral of register is
type arr is array(7 downto 0) of std_logic_vector(15 downto 0);
signal reg : arr : (others => '0');
begin


end Behavioral;

